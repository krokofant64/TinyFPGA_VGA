`include "K16Cpu.v"

`timescale 1 ns/10 ps  // time-unit = 1 ns, precision = 10 ps

module test2();

reg         clk;
reg         reset;
wire        hold;
wire        busy;
wire [15:0] address;
reg [15:0]  data_in;
wire [15:0] data_out;
wire        write;

always #1 clk = ~clk;

K16Cpu cpu(
  .clk(clk),
  .reset(reset),
  .hold(hold),
  .busy(busy),
  .address(address),
  .data_in(data_in),
  .data_out(data_out),
  .write(write));

  reg [15:0] ram[0:65535];

  always @(posedge clk)
    if (write) begin
      ram[address] <= data_out;
    end

  always @(posedge clk)
    data_in <= ram[address];

initial begin

//  ram[0]  = 16'hC38B;
//  ram[1]  = 16'hCB8B;
//  ram[2]  = 16'h6600;
//  ram[3]  = 16'h6E10;
//  ram[4]  = 16'h2900;
//  ram[5]  = 16'h4781;
//  ram[6]  = 16'h0480;
//  ram[7]  = 16'h2480;
//  ram[8]  = 16'h2903;
//  ram[9]  = 16'h0D8F;
//  ram[10] = 16'h4FFA;
//  ram[11] = 16'h9FFF;

//  ram[12] = 16'h002A;
//  ram[13] = 16'h00F3;

// ram[0] = 16'hC383;
// ram[1] = 16'h000C;
// ram[2] = 16'hE381;
// ram[3] = 16'h9FFF;
// ram[4] = 16'h000A;

ram[0] = 16'h7A10;
ram[1] = 16'hC386;
ram[2] = 16'hC786;
ram[3] = 16'hBC02;
ram[4] = 16'hEB85;
ram[5] = 16'h9FFF;
ram[6] = 16'h0810;
ram[7] = 16'h3C0D;
ram[8] = 16'h000A;
ram[9] = 16'h000D;


  $monitor("...clk=%b,reset=%b,hold=%b,busy=%b,address=%04X,data_in=%04X,data_out=%04X,write=%b,ram[9]=%04X,ram[10]=%04X,ram[16]=%04X",clk,reset,hold,busy,address,data_in,data_out,write,ram[9],ram[10],ram[16]);

  // initialize testbench variables
  clk = 1;
  reset = 1;

  #1
  clk = 0;
  reset = 0;

  repeat (50) @(posedge clk);
  $finish;

end
endmodule
