`ifndef SPRITE_V
`define SPRITE_V

module spriteBitmap(line, bits);
  input [3:0] line;
  output [63:0] bits;

  reg [63:0] rgbaBits[0:15]; // ROM array (64 x 16 bits)

  assign bits = rgbaBits[line];

  initial begin
    //                 RGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBA
    rgbaBits[0] <= 64'b0000000000000000000000000001000100010000000000000000000000000000;
    rgbaBits[1] <= 64'b0000000000000000000000011101110111010001000000000000000000000000;
    rgbaBits[2] <= 64'b0000000000000000000111011101110111011101000100000000000000000000;
    rgbaBits[3] <= 64'b0000000000000000000111010001110100011101000100000000000000000000;
    rgbaBits[4] <= 64'b0000000000000000000011011101110111011101000000000000000000000000;
    rgbaBits[5] <= 64'b0000000000000000000000001101000111010000000000000000000000000000;
    rgbaBits[6] <= 64'b0000000000001011101110111101110111011011101110110000000000000000;
    rgbaBits[7] <= 64'b0000000000001011000010111011101110111011000010110000000000000000;
    rgbaBits[8] <= 64'b0000000000001011000010111011111110111011000010110000000000000000;
    rgbaBits[9] <= 64'b0000000000001011000010111011111110111011000010110000000000000000;
    rgbaBits[10] <= 64'b0000000000001011000000110011010100110011000010110000000000000000;
    rgbaBits[11] <= 64'b0000000000001101000100010111011101110001000111010000000000000000;
    rgbaBits[12] <= 64'b0000000000000000000000010111000001110001000000000000000000000000;
    rgbaBits[13] <= 64'b0000000000000000000001110111000001110111000000000000000000000000;
    rgbaBits[14] <= 64'b0000000000000000000001110111000001110111000000000000000000000000;
    rgbaBits[15] <= 64'b0000000000000000000100010001000000010001000100000000000000000000;
    /*
    rgbaBits[0]    <= 64'b1101110111001100110011001100110010001000100010001000100010011001;
    rgbaBits[1]    <= 64'b1100110111011100110011001100110010001000100010001000100110011000;
    rgbaBits[2]    <= 64'b1100110011101110110011001100110010001000100010001001100110001000;
    rgbaBits[3]    <= 64'b1100110011001101110111001100110010001000100110011000100010001000;
    rgbaBits[4]    <= 64'b1100110011001100111111111111111110111011101110111000100010001000;
    rgbaBits[5]    <= 64'b1100110011001101111111111111111110111011101110111001100010001000;
    rgbaBits[6]    <= 64'b1100110011001101111111111111111110111011101110111001100010001000;
    rgbaBits[7]    <= 64'b1100110011011101111111111111111110111011101110111001100110001000;
    rgbaBits[8]    <= 64'b1000100010011001101110111011101100110011001100110001000100000000;
    rgbaBits[9]    <= 64'b1000100010001001101110111011101100110011001100110001000000000000;
    rgbaBits[10]   <= 64'b1000100010001001101110111011101100110011001100110000000000000000;
    rgbaBits[11]   <= 64'b1000100010001000101110111011101100110011001100110000000000000000;
    rgbaBits[12]   <= 64'b1000100010001000100110011000100000000000000000000001000100000000;
    rgbaBits[13]   <= 64'b1000100010011001100010001000100000000000000000000001000100000000;
    rgbaBits[14]   <= 64'b1000100110011000100010001000100000000000000000000000000100010000;
    rgbaBits[15]   <= 64'b1001100110001000100010001000100000000000000000000000000000010001;
    */
  end
endmodule

module drawSprite(line, column, red, green, blue, alpha);
  input [3:0] line;
  input [3:0] column;
  output red;
  output green;
  output blue;
  output alpha;

  wire [63:0] spriteBits;

  spriteBitmap bitmap(.line(line),
                      .bits(spriteBits));

  assign red   = spriteBits[{~column, 2'b00}];
  assign green = spriteBits[{~column, 2'b01}];
  assign blue  = spriteBits[{~column, 2'b10}];
  assign alpha = spriteBits[{~column, 2'b11}];

endmodule

module drawSprite2(line, column, red, green, blue, alpha);
  input [3:0] line;
  input [3:0] column;
  output red;
  output green;
  output blue;
  output alpha;

  reg [15:0] redbits[0:15]; // ROM array (16 x 16 bits)
  reg [15:0] greenbits[0:15]; // ROM array (16 x 16 bits)
  reg [15:0] bluebits[0:15]; // ROM array (16 x 16 bits)
  reg [15:0] alphabits[0:15]; // ROM array (16 x 16 bits)

  assign red    = redbits[line][~column];
  assign green  = greenbits[line][~column];
  assign blue   = bluebits[line][~column];
  assign alpha  = alphabits[line][~column];

  initial begin

    redbits[0]    <= 16'b1111111100000000;
    redbits[1]    <= 16'b1111111100000000;
    redbits[2]    <= 16'b1111111100000000;
    redbits[3]    <= 16'b1111111100000000;
    redbits[4]    <= 16'b1111111100000000;
    redbits[5]    <= 16'b1111111100000000;
    redbits[6]    <= 16'b1111111100000000;
    redbits[7]    <= 16'b1111111100000000;
    redbits[8]    <= 16'b1111111100000000;
    redbits[9]    <= 16'b1111111100000000;
    redbits[10]   <= 16'b1111111100000000;
    redbits[11]   <= 16'b1111111100000000;
    redbits[12]   <= 16'b1111111100000000;
    redbits[13]   <= 16'b1111111100000000;
    redbits[14]   <= 16'b1111111100000000;
    redbits[15]   <= 16'b1111111100000000;

    greenbits[0]  <= 16'b1111111111111111;
    greenbits[1]  <= 16'b1111111111111111;
    greenbits[2]  <= 16'b1111111111111111;
    greenbits[3]  <= 16'b1111111111111111;
    greenbits[4]  <= 16'b1111111111111111;
    greenbits[5]  <= 16'b1111111111111111;
    greenbits[6]  <= 16'b1111111111111111;
    greenbits[7]  <= 16'b1111111111111111;
    greenbits[8]  <= 16'b0000000000000000;
    greenbits[9]  <= 16'b0000000000000000;
    greenbits[10] <= 16'b0000000000000000;
    greenbits[11] <= 16'b0000000000000000;
    greenbits[12] <= 16'b0000000000000000;
    greenbits[13] <= 16'b0000000000000000;
    greenbits[14] <= 16'b0000000000000000;
    greenbits[15] <= 16'b0000000000000000;

    bluebits[0]   <= 16'b0000000000000000;
    bluebits[1]   <= 16'b0000000000000000;
    bluebits[2]   <= 16'b0000000000000000;
    bluebits[3]   <= 16'b0000000000000000;
    bluebits[4]   <= 16'b0000111111110000;
    bluebits[5]   <= 16'b0000111111110000;
    bluebits[6]   <= 16'b0000111111110000;
    bluebits[7]   <= 16'b0000111111110000;
    bluebits[8]   <= 16'b0000111111110000;
    bluebits[9]   <= 16'b0000111111110000;
    bluebits[10]  <= 16'b0000111111110000;
    bluebits[11]  <= 16'b0000111111110000;
    bluebits[12]  <= 16'b0000000000000000;
    bluebits[13]  <= 16'b0000000000000000;
    bluebits[14]  <= 16'b0000000000000000;
    bluebits[15]  <= 16'b0000000000000000;

    alphabits[0]  <= 16'b1100000000000011;
    alphabits[1]  <= 16'b0110000000000110;
    alphabits[2]  <= 16'b0011000000001100;
    alphabits[3]  <= 16'b0001100000110000;
    alphabits[4]  <= 16'b0000111111110000;
    alphabits[5]  <= 16'b0001111111111000;
    alphabits[6]  <= 16'b0001111111111000;
    alphabits[7]  <= 16'b0011111111111100;
    alphabits[8]  <= 16'b0011111111111100;
    alphabits[9]  <= 16'b0001111111111000;
    alphabits[10] <= 16'b0001111111111000;
    alphabits[11] <= 16'b0000111111110000;
    alphabits[12] <= 16'b0001100000011000;
    alphabits[13] <= 16'b0011000000001100;
    alphabits[14] <= 16'b0110000000000110;
    alphabits[15] <= 16'b1100000000000011;

  end
endmodule

`endif
