`ifndef SPRITE_V
`define SPRITE_V

module SpriteBitmap(line, bits);
  input [3:0] line;
  output [63:0] bits;

  reg [63:0] rgbaBits[0:15]; // ROM array (64 x 16 bits)

  assign bits = rgbaBits[line];

  initial begin
    //                 RGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBARGBA
    rgbaBits[0] <= 64'b0000000000000000000000000001000100010000000000000000000000000000;
    rgbaBits[1] <= 64'b0000000000000000000000011101110111010001000000000000000000000000;
    rgbaBits[2] <= 64'b0000000000000000000111011101110111011101000100000000000000000000;
    rgbaBits[3] <= 64'b0000000000000000000111010001110100011101000100000000000000000000;
    rgbaBits[4] <= 64'b0000000000000000000011011101110111011101000000000000000000000000;
    rgbaBits[5] <= 64'b0000000000000000000000001101000111010000000000000000000000000000;
    rgbaBits[6] <= 64'b0000000000001011101110111101110111011011101110110000000000000000;
    rgbaBits[7] <= 64'b0000000000001011000010111011101110111011000010110000000000000000;
    rgbaBits[8] <= 64'b0000000000001011000010111011111110111011000010110000000000000000;
    rgbaBits[9] <= 64'b0000000000001011000010111011111110111011000010110000000000000000;
    rgbaBits[10] <= 64'b0000000000001011000000110011010100110011000010110000000000000000;
    rgbaBits[11] <= 64'b0000000000001101000100010111011101110001000111010000000000000000;
    rgbaBits[12] <= 64'b0000000000000000000000010111000001110001000000000000000000000000;
    rgbaBits[13] <= 64'b0000000000000000000001110111000001110111000000000000000000000000;
    rgbaBits[14] <= 64'b0000000000000000000001110111000001110111000000000000000000000000;
    rgbaBits[15] <= 64'b0000000000000000000100010001000000010001000100000000000000000000;
  end
endmodule
`endif
